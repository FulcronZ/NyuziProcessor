// 
// Copyright 2015 Pipat Methavanitpong
// 
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     http://www.apache.org/licenses/LICENSE-2.0
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 

/// An asynchronous counter

module counter
	#(parameter WIDTH = 32)
	(input						reset,
	input						increment,
	input						enable,
	output logic[WIDTH - 1:0] 	value);
	
	always_ff @(posedge increment, posedge reset)
	begin : update
		if (reset)
			value <= 0;
		else
			if (enable)
				value <= value + 1;
		end
	end
endmodule
